// (C) 2001-2012 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License Subscription 
// Agreement, Altera MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


// $Id: //acds/rel/12.1/ip/merlin/altera_merlin_router/altera_merlin_router.sv.terp#1 $
// $Revision: #1 $
// $Date: 2012/08/12 $
// $Author: swbranch $

// -------------------------------------------------------
// Merlin Router
//
// Asserts the appropriate one-hot encoded channel based on 
// either (a) the address or (b) the dest id. The DECODER_TYPE
// parameter controls this behaviour. 0 means address decoder,
// 1 means dest id decoder.
//
// In the case of (a), it also sets the destination id.
// -------------------------------------------------------

`timescale 1 ns / 1 ns

module first_nios2_system_addr_router_001_default_decode
  #(
     parameter DEFAULT_CHANNEL = 1,
               DEFAULT_DESTID = 1 
   )
<<<<<<< HEAD
  (output [87 - 85 : 0] default_destination_id,
   output [6-1 : 0] default_src_channel
=======
  (output [85 - 83 : 0] default_destination_id,
   output [7-1 : 0] default_src_channel
>>>>>>> 5f0fa4d91aa97f188f2e619db808c790c0793725
  );

  assign default_destination_id = 
    DEFAULT_DESTID[87 - 85 : 0];
  generate begin : default_decode
    if (DEFAULT_CHANNEL == -1)
      assign default_src_channel = '0;
    else
<<<<<<< HEAD
      assign default_src_channel = 6'b1 << DEFAULT_CHANNEL;
  end
  endgenerate
=======
      assign default_src_channel = 7'b1 << DEFAULT_CHANNEL;
  end endgenerate
>>>>>>> 5f0fa4d91aa97f188f2e619db808c790c0793725

endmodule


module first_nios2_system_addr_router_001
(
    // -------------------
    // Clock & Reset
    // -------------------
    input clk,
    input reset,

    // -------------------
    // Command Sink (Input)
    // -------------------
    input                       sink_valid,
    input  [98-1 : 0]    sink_data,
    input                       sink_startofpacket,
    input                       sink_endofpacket,
    output                      sink_ready,

    // -------------------
    // Command Source (Output)
    // -------------------
    output                          src_valid,
<<<<<<< HEAD
    output reg [98-1    : 0] src_data,
    output reg [6-1 : 0] src_channel,
=======
    output reg [96-1    : 0] src_data,
    output reg [7-1 : 0] src_channel,
>>>>>>> 5f0fa4d91aa97f188f2e619db808c790c0793725
    output                          src_startofpacket,
    output                          src_endofpacket,
    input                           src_ready
);

    // -------------------------------------------------------
    // Local parameters and variables
    // -------------------------------------------------------
    localparam PKT_ADDR_H = 60;
    localparam PKT_ADDR_L = 36;
<<<<<<< HEAD
    localparam PKT_DEST_ID_H = 87;
    localparam PKT_DEST_ID_L = 85;
    localparam ST_DATA_W = 98;
    localparam ST_CHANNEL_W = 6;
=======
    localparam PKT_DEST_ID_H = 85;
    localparam PKT_DEST_ID_L = 83;
    localparam ST_DATA_W = 96;
    localparam ST_CHANNEL_W = 7;
>>>>>>> 5f0fa4d91aa97f188f2e619db808c790c0793725
    localparam DECODER_TYPE = 0;

    localparam PKT_TRANS_WRITE = 63;
    localparam PKT_TRANS_READ  = 64;

    localparam PKT_ADDR_W = PKT_ADDR_H-PKT_ADDR_L + 1;
    localparam PKT_DEST_ID_W = PKT_DEST_ID_H-PKT_DEST_ID_L + 1;




    // -------------------------------------------------------
    // Figure out the number of bits to mask off for each slave span
    // during address decoding
    // -------------------------------------------------------
<<<<<<< HEAD
    localparam PAD0 = log2ceil(64'h1000000 - 64'h800000);
    localparam PAD1 = log2ceil(64'h1001000 - 64'h1000800);
    localparam PAD2 = log2ceil(64'h1001020 - 64'h1001000);
    localparam PAD3 = log2ceil(64'h1001030 - 64'h1001020);
    localparam PAD4 = log2ceil(64'h1001038 - 64'h1001030);
    localparam PAD5 = log2ceil(64'h1001040 - 64'h1001038);
=======
    localparam PAD0 = log2ceil(32'h10 - 32'h0);
    localparam PAD1 = log2ceil(32'h1000000 - 32'h800000);
    localparam PAD2 = log2ceil(32'h1001000 - 32'h1000800);
    localparam PAD3 = log2ceil(32'h1001020 - 32'h1001000);
    localparam PAD4 = log2ceil(32'h1001030 - 32'h1001020);
    localparam PAD5 = log2ceil(32'h1001038 - 32'h1001030);
    localparam PAD6 = log2ceil(32'h1001040 - 32'h1001038);

>>>>>>> 5f0fa4d91aa97f188f2e619db808c790c0793725
    // -------------------------------------------------------
    // Work out which address bits are significant based on the
    // address range of the slaves. If the required width is too
    // large or too small, we use the address field width instead.
    // -------------------------------------------------------
    localparam ADDR_RANGE = 64'h1001040;
    localparam RANGE_ADDR_WIDTH = log2ceil(ADDR_RANGE);
    localparam OPTIMIZED_ADDR_H = (RANGE_ADDR_WIDTH > PKT_ADDR_W) ||
                                  (RANGE_ADDR_WIDTH == 0) ?
                                        PKT_ADDR_H :
                                        PKT_ADDR_L + RANGE_ADDR_WIDTH - 1;
    localparam RG = RANGE_ADDR_WIDTH-1;

      wire [PKT_ADDR_W-1 : 0] address = sink_data[OPTIMIZED_ADDR_H : PKT_ADDR_L];

    // -------------------------------------------------------
    // Pass almost everything through, untouched
    // -------------------------------------------------------
    assign sink_ready        = src_ready;
    assign src_valid         = sink_valid;
    assign src_startofpacket = sink_startofpacket;
    assign src_endofpacket   = sink_endofpacket;

    wire [PKT_DEST_ID_W-1:0] default_destid;
    wire [7-1 : 0] default_src_channel;




    first_nios2_system_addr_router_001_default_decode the_default_decode(
      .default_destination_id (default_destid),
      .default_src_channel (default_src_channel)
    );

    always @* begin
        src_data    = sink_data;
        src_channel = default_src_channel;

        src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = default_destid;
        // --------------------------------------------------
        // Address Decoder
        // Sets the channel and destination ID based on the address
        // --------------------------------------------------

        // ( 0x0 .. 0x10 )
        if ( {address[RG:PAD0],{PAD0{1'b0}}} == 'h0 ) begin
            src_channel = 7'b1000000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 6;
        end

        // ( 0x800000 .. 0x1000000 )
<<<<<<< HEAD
        if ( {address[RG:PAD0],{PAD0{1'b0}}} == 25'h800000 ) begin
            src_channel = 6'b000010;
=======
        if ( {address[RG:PAD1],{PAD1{1'b0}}} == 'h800000 ) begin
            src_channel = 7'b0000010;
>>>>>>> 5f0fa4d91aa97f188f2e619db808c790c0793725
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 1;
        end

        // ( 0x1000800 .. 0x1001000 )
<<<<<<< HEAD
        if ( {address[RG:PAD1],{PAD1{1'b0}}} == 25'h1000800 ) begin
            src_channel = 6'b000001;
=======
        if ( {address[RG:PAD2],{PAD2{1'b0}}} == 'h1000800 ) begin
            src_channel = 7'b0000001;
>>>>>>> 5f0fa4d91aa97f188f2e619db808c790c0793725
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 0;
        end

        // ( 0x1001000 .. 0x1001020 )
<<<<<<< HEAD
        if ( {address[RG:PAD2],{PAD2{1'b0}}} == 25'h1001000 ) begin
            src_channel = 6'b010000;
=======
        if ( {address[RG:PAD3],{PAD3{1'b0}}} == 'h1001000 ) begin
            src_channel = 7'b0010000;
>>>>>>> 5f0fa4d91aa97f188f2e619db808c790c0793725
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 4;
        end

        // ( 0x1001020 .. 0x1001030 )
<<<<<<< HEAD
        if ( {address[RG:PAD3],{PAD3{1'b0}}} == 25'h1001020 ) begin
            src_channel = 6'b100000;
=======
        if ( {address[RG:PAD4],{PAD4{1'b0}}} == 'h1001020 ) begin
            src_channel = 7'b0100000;
>>>>>>> 5f0fa4d91aa97f188f2e619db808c790c0793725
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 5;
        end

        // ( 0x1001030 .. 0x1001038 )
<<<<<<< HEAD
        if ( {address[RG:PAD4],{PAD4{1'b0}}} == 25'h1001030 ) begin
            src_channel = 6'b000100;
=======
        if ( {address[RG:PAD5],{PAD5{1'b0}}} == 'h1001030 ) begin
            src_channel = 7'b0000100;
>>>>>>> 5f0fa4d91aa97f188f2e619db808c790c0793725
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 2;
        end

        // ( 0x1001038 .. 0x1001040 )
<<<<<<< HEAD
        if ( {address[RG:PAD5],{PAD5{1'b0}}} == 25'h1001038 ) begin
            src_channel = 6'b001000;
=======
        if ( {address[RG:PAD6],{PAD6{1'b0}}} == 'h1001038 ) begin
            src_channel = 7'b0001000;
>>>>>>> 5f0fa4d91aa97f188f2e619db808c790c0793725
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 3;
        end

end


    // --------------------------------------------------
    // Ceil(log2()) function
    // --------------------------------------------------
    function integer log2ceil;
        input reg[65:0] val;
        reg [65:0] i;

        begin
            i = 1;
            log2ceil = 0;

            while (i < val) begin
                log2ceil = log2ceil + 1;
                i = i << 1;
            end
        end
    endfunction

endmodule


